library verilog;
use verilog.vl_types.all;
entity DECODER2_4_vlg_vec_tst is
end DECODER2_4_vlg_vec_tst;
