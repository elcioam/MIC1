library verilog;
use verilog.vl_types.all;
entity REGISTER_32BIT_vlg_vec_tst is
end REGISTER_32BIT_vlg_vec_tst;
